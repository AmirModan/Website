-- internal_pin_if.vhd

-- Generated using ACDS version 19.1 670

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity internal_pin_if is
	port (
		clk_clk                      : in  std_logic                     := '0';             --                   clk.clk
		led31_to_0_export            : in  std_logic_vector(31 downto 0) := (others => '0'); --            led31_to_0.export
		led63_to_32_export           : in  std_logic_vector(31 downto 0) := (others => '0'); --           led63_to_32.export
		param1_export                : out std_logic_vector(31 downto 0);                    --                param1.export
		param2_export                : out std_logic_vector(31 downto 0);                    --                param2.export
		param3_export                : out std_logic_vector(31 downto 0);                    --                param3.export
		pbs11_to_10_sws9_to_0_export : out std_logic_vector(11 downto 0);                    -- pbs11_to_10_sws9_to_0.export
		reset_reset_n                : in  std_logic                     := '0'              --                 reset.reset_n
	);
end entity internal_pin_if;

architecture rtl of internal_pin_if is
	component internal_pin_if_JTAG_2_Avalon_IP is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component internal_pin_if_JTAG_2_Avalon_IP;

	component internal_pin_if_LED_IP_0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component internal_pin_if_LED_IP_0;

	component internal_pin_if_SW_IP is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(11 downto 0)                     -- export
		);
	end component internal_pin_if_SW_IP;

	component internal_pin_if_param1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component internal_pin_if_param1;

	component internal_pin_if_mm_interconnect_0 is
		port (
			CLK_IP_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			JTAG_2_Avalon_IP_clk_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			JTAG_2_Avalon_IP_master_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			LED_IP_0_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			JTAG_2_Avalon_IP_master_address                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			JTAG_2_Avalon_IP_master_waitrequest                                  : out std_logic;                                        -- waitrequest
			JTAG_2_Avalon_IP_master_byteenable                                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			JTAG_2_Avalon_IP_master_read                                         : in  std_logic                     := 'X';             -- read
			JTAG_2_Avalon_IP_master_readdata                                     : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_2_Avalon_IP_master_readdatavalid                                : out std_logic;                                        -- readdatavalid
			JTAG_2_Avalon_IP_master_write                                        : in  std_logic                     := 'X';             -- write
			JTAG_2_Avalon_IP_master_writedata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			LED_IP_0_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			LED_IP_0_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LED_IP_1_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			LED_IP_1_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			param1_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			param1_s1_write                                                      : out std_logic;                                        -- write
			param1_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			param1_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			param1_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			param2_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			param2_s1_write                                                      : out std_logic;                                        -- write
			param2_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			param2_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			param2_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			param3_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			param3_s1_write                                                      : out std_logic;                                        -- write
			param3_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			param3_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			param3_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			SW_IP_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			SW_IP_s1_write                                                       : out std_logic;                                        -- write
			SW_IP_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SW_IP_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			SW_IP_s1_chipselect                                                  : out std_logic                                         -- chipselect
		);
	end component internal_pin_if_mm_interconnect_0;

	component internal_pin_if_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component internal_pin_if_rst_controller;

	component internal_pin_if_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component internal_pin_if_rst_controller_001;

	signal jtag_2_avalon_ip_master_readdata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_2_Avalon_IP_master_readdata -> JTAG_2_Avalon_IP:master_readdata
	signal jtag_2_avalon_ip_master_waitrequest          : std_logic;                     -- mm_interconnect_0:JTAG_2_Avalon_IP_master_waitrequest -> JTAG_2_Avalon_IP:master_waitrequest
	signal jtag_2_avalon_ip_master_address              : std_logic_vector(31 downto 0); -- JTAG_2_Avalon_IP:master_address -> mm_interconnect_0:JTAG_2_Avalon_IP_master_address
	signal jtag_2_avalon_ip_master_read                 : std_logic;                     -- JTAG_2_Avalon_IP:master_read -> mm_interconnect_0:JTAG_2_Avalon_IP_master_read
	signal jtag_2_avalon_ip_master_byteenable           : std_logic_vector(3 downto 0);  -- JTAG_2_Avalon_IP:master_byteenable -> mm_interconnect_0:JTAG_2_Avalon_IP_master_byteenable
	signal jtag_2_avalon_ip_master_readdatavalid        : std_logic;                     -- mm_interconnect_0:JTAG_2_Avalon_IP_master_readdatavalid -> JTAG_2_Avalon_IP:master_readdatavalid
	signal jtag_2_avalon_ip_master_write                : std_logic;                     -- JTAG_2_Avalon_IP:master_write -> mm_interconnect_0:JTAG_2_Avalon_IP_master_write
	signal jtag_2_avalon_ip_master_writedata            : std_logic_vector(31 downto 0); -- JTAG_2_Avalon_IP:master_writedata -> mm_interconnect_0:JTAG_2_Avalon_IP_master_writedata
	signal mm_interconnect_0_led_ip_0_s1_readdata       : std_logic_vector(31 downto 0); -- LED_IP_0:readdata -> mm_interconnect_0:LED_IP_0_s1_readdata
	signal mm_interconnect_0_led_ip_0_s1_address        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LED_IP_0_s1_address -> LED_IP_0:address
	signal mm_interconnect_0_sw_ip_s1_chipselect        : std_logic;                     -- mm_interconnect_0:SW_IP_s1_chipselect -> SW_IP:chipselect
	signal mm_interconnect_0_sw_ip_s1_readdata          : std_logic_vector(31 downto 0); -- SW_IP:readdata -> mm_interconnect_0:SW_IP_s1_readdata
	signal mm_interconnect_0_sw_ip_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SW_IP_s1_address -> SW_IP:address
	signal mm_interconnect_0_sw_ip_s1_write             : std_logic;                     -- mm_interconnect_0:SW_IP_s1_write -> mm_interconnect_0_sw_ip_s1_write:in
	signal mm_interconnect_0_sw_ip_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:SW_IP_s1_writedata -> SW_IP:writedata
	signal mm_interconnect_0_led_ip_1_s1_readdata       : std_logic_vector(31 downto 0); -- LED_IP_1:readdata -> mm_interconnect_0:LED_IP_1_s1_readdata
	signal mm_interconnect_0_led_ip_1_s1_address        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LED_IP_1_s1_address -> LED_IP_1:address
	signal mm_interconnect_0_param1_s1_chipselect       : std_logic;                     -- mm_interconnect_0:param1_s1_chipselect -> param1:chipselect
	signal mm_interconnect_0_param1_s1_readdata         : std_logic_vector(31 downto 0); -- param1:readdata -> mm_interconnect_0:param1_s1_readdata
	signal mm_interconnect_0_param1_s1_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:param1_s1_address -> param1:address
	signal mm_interconnect_0_param1_s1_write            : std_logic;                     -- mm_interconnect_0:param1_s1_write -> mm_interconnect_0_param1_s1_write:in
	signal mm_interconnect_0_param1_s1_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:param1_s1_writedata -> param1:writedata
	signal mm_interconnect_0_param2_s1_chipselect       : std_logic;                     -- mm_interconnect_0:param2_s1_chipselect -> param2:chipselect
	signal mm_interconnect_0_param2_s1_readdata         : std_logic_vector(31 downto 0); -- param2:readdata -> mm_interconnect_0:param2_s1_readdata
	signal mm_interconnect_0_param2_s1_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:param2_s1_address -> param2:address
	signal mm_interconnect_0_param2_s1_write            : std_logic;                     -- mm_interconnect_0:param2_s1_write -> mm_interconnect_0_param2_s1_write:in
	signal mm_interconnect_0_param2_s1_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:param2_s1_writedata -> param2:writedata
	signal mm_interconnect_0_param3_s1_chipselect       : std_logic;                     -- mm_interconnect_0:param3_s1_chipselect -> param3:chipselect
	signal mm_interconnect_0_param3_s1_readdata         : std_logic_vector(31 downto 0); -- param3:readdata -> mm_interconnect_0:param3_s1_readdata
	signal mm_interconnect_0_param3_s1_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:param3_s1_address -> param3:address
	signal mm_interconnect_0_param3_s1_write            : std_logic;                     -- mm_interconnect_0:param3_s1_write -> mm_interconnect_0_param3_s1_write:in
	signal mm_interconnect_0_param3_s1_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:param3_s1_writedata -> param3:writedata
	signal rst_controller_reset_out_reset               : std_logic;                     -- rst_controller:reset_out -> JTAG_2_Avalon_IP:clk_reset_reset
	signal jtag_2_avalon_ip_master_reset_reset          : std_logic;                     -- JTAG_2_Avalon_IP:master_reset_reset -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset           : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:LED_IP_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset           : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:JTAG_2_Avalon_IP_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:JTAG_2_Avalon_IP_master_translator_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                      : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_sw_ip_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_sw_ip_s1_write:inv -> SW_IP:write_n
	signal mm_interconnect_0_param1_s1_write_ports_inv  : std_logic;                     -- mm_interconnect_0_param1_s1_write:inv -> param1:write_n
	signal mm_interconnect_0_param2_s1_write_ports_inv  : std_logic;                     -- mm_interconnect_0_param2_s1_write:inv -> param2:write_n
	signal mm_interconnect_0_param3_s1_write_ports_inv  : std_logic;                     -- mm_interconnect_0_param3_s1_write:inv -> param3:write_n
	signal rst_controller_001_reset_out_reset_ports_inv : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [LED_IP_0:reset_n, LED_IP_1:reset_n, SW_IP:reset_n, param1:reset_n, param2:reset_n, param3:reset_n]

begin

	jtag_2_avalon_ip : component internal_pin_if_JTAG_2_Avalon_IP
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                               --          clk.clk
			clk_reset_reset      => rst_controller_reset_out_reset,        --    clk_reset.reset
			master_address       => jtag_2_avalon_ip_master_address,       --       master.address
			master_readdata      => jtag_2_avalon_ip_master_readdata,      --             .readdata
			master_read          => jtag_2_avalon_ip_master_read,          --             .read
			master_write         => jtag_2_avalon_ip_master_write,         --             .write
			master_writedata     => jtag_2_avalon_ip_master_writedata,     --             .writedata
			master_waitrequest   => jtag_2_avalon_ip_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_2_avalon_ip_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_2_avalon_ip_master_byteenable,    --             .byteenable
			master_reset_reset   => jtag_2_avalon_ip_master_reset_reset    -- master_reset.reset
		);

	led_ip_0 : component internal_pin_if_LED_IP_0
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_led_ip_0_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_led_ip_0_s1_readdata,       --                    .readdata
			in_port  => led31_to_0_export                             -- external_connection.export
		);

	led_ip_1 : component internal_pin_if_LED_IP_0
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_led_ip_1_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_led_ip_1_s1_readdata,       --                    .readdata
			in_port  => led63_to_32_export                            -- external_connection.export
		);

	sw_ip : component internal_pin_if_SW_IP
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_sw_ip_s1_address,           --                  s1.address
			write_n    => mm_interconnect_0_sw_ip_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_0_sw_ip_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_0_sw_ip_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_0_sw_ip_s1_readdata,          --                    .readdata
			out_port   => pbs11_to_10_sws9_to_0_export                  -- external_connection.export
		);

	param1 : component internal_pin_if_param1
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_param1_s1_address,          --                  s1.address
			write_n    => mm_interconnect_0_param1_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_0_param1_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_0_param1_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_0_param1_s1_readdata,         --                    .readdata
			out_port   => param1_export                                 -- external_connection.export
		);

	param2 : component internal_pin_if_param1
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_param2_s1_address,          --                  s1.address
			write_n    => mm_interconnect_0_param2_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_0_param2_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_0_param2_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_0_param2_s1_readdata,         --                    .readdata
			out_port   => param2_export                                 -- external_connection.export
		);

	param3 : component internal_pin_if_param1
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_param3_s1_address,          --                  s1.address
			write_n    => mm_interconnect_0_param3_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_0_param3_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_0_param3_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_0_param3_s1_readdata,         --                    .readdata
			out_port   => param3_export                                 -- external_connection.export
		);

	mm_interconnect_0 : component internal_pin_if_mm_interconnect_0
		port map (
			CLK_IP_clk_clk                                                       => clk_clk,                                --                                                     CLK_IP_clk.clk
			JTAG_2_Avalon_IP_clk_reset_reset_bridge_in_reset_reset               => rst_controller_002_reset_out_reset,     --               JTAG_2_Avalon_IP_clk_reset_reset_bridge_in_reset.reset
			JTAG_2_Avalon_IP_master_translator_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,     -- JTAG_2_Avalon_IP_master_translator_reset_reset_bridge_in_reset.reset
			LED_IP_0_reset_reset_bridge_in_reset_reset                           => rst_controller_001_reset_out_reset,     --                           LED_IP_0_reset_reset_bridge_in_reset.reset
			JTAG_2_Avalon_IP_master_address                                      => jtag_2_avalon_ip_master_address,        --                                        JTAG_2_Avalon_IP_master.address
			JTAG_2_Avalon_IP_master_waitrequest                                  => jtag_2_avalon_ip_master_waitrequest,    --                                                               .waitrequest
			JTAG_2_Avalon_IP_master_byteenable                                   => jtag_2_avalon_ip_master_byteenable,     --                                                               .byteenable
			JTAG_2_Avalon_IP_master_read                                         => jtag_2_avalon_ip_master_read,           --                                                               .read
			JTAG_2_Avalon_IP_master_readdata                                     => jtag_2_avalon_ip_master_readdata,       --                                                               .readdata
			JTAG_2_Avalon_IP_master_readdatavalid                                => jtag_2_avalon_ip_master_readdatavalid,  --                                                               .readdatavalid
			JTAG_2_Avalon_IP_master_write                                        => jtag_2_avalon_ip_master_write,          --                                                               .write
			JTAG_2_Avalon_IP_master_writedata                                    => jtag_2_avalon_ip_master_writedata,      --                                                               .writedata
			LED_IP_0_s1_address                                                  => mm_interconnect_0_led_ip_0_s1_address,  --                                                    LED_IP_0_s1.address
			LED_IP_0_s1_readdata                                                 => mm_interconnect_0_led_ip_0_s1_readdata, --                                                               .readdata
			LED_IP_1_s1_address                                                  => mm_interconnect_0_led_ip_1_s1_address,  --                                                    LED_IP_1_s1.address
			LED_IP_1_s1_readdata                                                 => mm_interconnect_0_led_ip_1_s1_readdata, --                                                               .readdata
			param1_s1_address                                                    => mm_interconnect_0_param1_s1_address,    --                                                      param1_s1.address
			param1_s1_write                                                      => mm_interconnect_0_param1_s1_write,      --                                                               .write
			param1_s1_readdata                                                   => mm_interconnect_0_param1_s1_readdata,   --                                                               .readdata
			param1_s1_writedata                                                  => mm_interconnect_0_param1_s1_writedata,  --                                                               .writedata
			param1_s1_chipselect                                                 => mm_interconnect_0_param1_s1_chipselect, --                                                               .chipselect
			param2_s1_address                                                    => mm_interconnect_0_param2_s1_address,    --                                                      param2_s1.address
			param2_s1_write                                                      => mm_interconnect_0_param2_s1_write,      --                                                               .write
			param2_s1_readdata                                                   => mm_interconnect_0_param2_s1_readdata,   --                                                               .readdata
			param2_s1_writedata                                                  => mm_interconnect_0_param2_s1_writedata,  --                                                               .writedata
			param2_s1_chipselect                                                 => mm_interconnect_0_param2_s1_chipselect, --                                                               .chipselect
			param3_s1_address                                                    => mm_interconnect_0_param3_s1_address,    --                                                      param3_s1.address
			param3_s1_write                                                      => mm_interconnect_0_param3_s1_write,      --                                                               .write
			param3_s1_readdata                                                   => mm_interconnect_0_param3_s1_readdata,   --                                                               .readdata
			param3_s1_writedata                                                  => mm_interconnect_0_param3_s1_writedata,  --                                                               .writedata
			param3_s1_chipselect                                                 => mm_interconnect_0_param3_s1_chipselect, --                                                               .chipselect
			SW_IP_s1_address                                                     => mm_interconnect_0_sw_ip_s1_address,     --                                                       SW_IP_s1.address
			SW_IP_s1_write                                                       => mm_interconnect_0_sw_ip_s1_write,       --                                                               .write
			SW_IP_s1_readdata                                                    => mm_interconnect_0_sw_ip_s1_readdata,    --                                                               .readdata
			SW_IP_s1_writedata                                                   => mm_interconnect_0_sw_ip_s1_writedata,   --                                                               .writedata
			SW_IP_s1_chipselect                                                  => mm_interconnect_0_sw_ip_s1_chipselect   --                                                               .chipselect
		);

	rst_controller : component internal_pin_if_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => jtag_2_avalon_ip_master_reset_reset, -- reset_in1.reset
			clk            => open,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_001 : component internal_pin_if_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component internal_pin_if_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => jtag_2_avalon_ip_master_reset_reset, -- reset_in1.reset
			clk            => clk_clk,                             --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_sw_ip_s1_write_ports_inv <= not mm_interconnect_0_sw_ip_s1_write;

	mm_interconnect_0_param1_s1_write_ports_inv <= not mm_interconnect_0_param1_s1_write;

	mm_interconnect_0_param2_s1_write_ports_inv <= not mm_interconnect_0_param2_s1_write;

	mm_interconnect_0_param3_s1_write_ports_inv <= not mm_interconnect_0_param3_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of internal_pin_if
